class transmit_dynamic_frame_test extends uart_base_test;
	`uvm_component_utils(transmit_dynamic_frame_test)
	
	uvm_status_e       status;
	uart_configuration uart_config2;
	vip_tx_sequence		 seq;

	//----------------------------------------
	// Constructor
	//----------------------------------------
	function new(string name = "transmit_dynamic_frame_test", uvm_component parent);
		super.new(name,parent);
	endfunction

	//-------------------------------------
	// run phase
	//-------------------------------------
	virtual task run_phase(uvm_phase phase);
		bit[7:0]  transmit_data;
		bit[5:0]  transmit_data2;
		bit[4:0]  transmit_data3;
		bit[31:0] rdata;
		phase.raise_objection(this);
		
		// config VIP
		uart_config2 = uart_configuration::type_id::create("uart_config2");
		uart_config2.baud_rate   = 115200;
		uart_config2.data_width  = 8;
		uart_config2.parity_mode = uart_configuration::PARITY_NONE;
		uart_config2.stop_bits   = 1;
		`uvm_info(get_type_name(),"UART agent updating...",UVM_LOW)
		env.uart_agt.update_config(uart_config2);
		// config DUT
		regmodel.MDR.write(status,32'h00); #50ns;
		regmodel.DLL.write(status,32'h36); #50ns;
		regmodel.LCR.write(status,32'h33); #50ns;
	
		transmit_data = $urandom();
		regmodel.TBR.write(status,transmit_data);
			
		#((1.0e9/uart_config2.baud_rate)*13ns);

		// reconfig VIP to change frame
		uart_config2.data_width = 6;
		uart_config2.stop_bits  = 2;
		`uvm_info(get_type_name(),"UART agent updating...",UVM_LOW)
		env.uart_agt.update_config(uart_config2);
		// reconfig DUT to change frame
		transmit_data2 = $urandom();
		regmodel.LCR.write(status,32'h25);
		regmodel.TBR.write(status,transmit_data2);

		#((1.0e9/uart_config2.baud_rate)*13ns);

		// reconfig VIP to change frame
		uart_config2.data_width = 5;
		uart_config2.stop_bits  = 1;
		`uvm_info(get_type_name(),"UART agent updating...",UVM_LOW)
		env.uart_agt.update_config(uart_config2);
		// reconfig DUT to change frame
		transmit_data3 = $urandom();
		regmodel.LCR.write(status,32'h20);
		regmodel.TBR.write(status,transmit_data3);

		#((1.0e9/uart_config2.baud_rate)*13ns);

		phase.drop_objection(this);
	endtask

endclass
