class dis_rx_fifo_full_interrupt_test extends uart_base_test;
	`uvm_component_utils(dis_rx_fifo_full_interrupt_test)
	
	uvm_status_e       status;
	uart_configuration uart_config2;
	vip_tx_sequence		 seq;

	//----------------------------------------
	// Constructor
	//----------------------------------------
	function new(string name = "dis_rx_fifo_full_interrupt_test", uvm_component parent);
		super.new(name,parent);
	endfunction

	//-------------------------------------
	// run phase
	//-------------------------------------
	virtual task run_phase(uvm_phase phase);
		bit[7:0] rdata;
		phase.raise_objection(this);

		wait(ahb_vif.HRESETn === 1);

		// config VIP
		uart_config2 = uart_configuration::type_id::create("uart_config2");
		uart_config2.baud_rate   = 115200;
		uart_config2.data_width  = 8;
		uart_config2.parity_mode = uart_configuration::PARITY_EVEN;
		uart_config2.stop_bits   = 2;
		`uvm_info(get_type_name(),"UART agent updating...",UVM_LOW)
		env.uart_agt.update_config(uart_config2);
		// config DUT
		regmodel.IER.write(status,32'h00); #1ns;
		if(uart_vif.interrupt === 0) // check before rx fifo not full
			`uvm_info(get_type_name(),"RX FIFO is not full, interrupt is disable so interrupt = 0",UVM_LOW)
		else
			`uvm_error(get_type_name(),"RX FIFO is not full, interrupt must equal 0")
		regmodel.FSR.read(status,rdata);
		if(rdata[2] === 0)
			`uvm_info(get_type_name(),"RX FIFO is not full, rx fifo full status = 0",UVM_LOW)
		else
			`uvm_error(get_type_name(),"RX FIFO is not full, rx fifo full status must equal 0")

		regmodel.MDR.write(status,32'h00); #(50*1ns);
		regmodel.DLL.write(status,32'h36); #(50*1ns);
		regmodel.LCR.write(status,32'h3F); #(50*1ns);

		seq = vip_tx_sequence::type_id::create("seq");
		
		repeat(16) seq.start(env.uart_agt.uart_seqcer);

		if(uart_vif.interrupt === 1) // check rx fifo full
			`uvm_error(get_type_name(),"RX FIFO full but interrupt is disable, interrupt cannot trigger")
		regmodel.FSR.read(status,rdata);
		if(rdata[2] === 1)
			`uvm_info(get_type_name(),"RX FIFO has data, rx fifo full status trigger to 1",UVM_LOW)
		else
			`uvm_error(get_type_name(),"RX FIFO has data, rx fifo full status must be = 1")
		
		regmodel.RBR.read(status,rdata);
		env.uart_sb.update_rbr_data(rdata);

		#1ns;
		if(uart_vif.interrupt === 0) // check rx fifo not full
			`uvm_info(get_type_name(),"RX FIFO is not full, interrupt is disable so interrupt = 0",UVM_LOW)
		else
			`uvm_error(get_type_name(),"RX FIFO is not full, interrupt is disable so interrupt must equal 0")
		regmodel.FSR.read(status,rdata);
		if(rdata[2] === 0)
			`uvm_info(get_type_name(),"RX FIFO is not full, rx fifo full status = 0",UVM_LOW)
		else
			`uvm_error(get_type_name(),"RX FIFO is not full, rx fifo full status must equal 0")

		repeat(15) begin
			regmodel.RBR.read(status,rdata);
			env.uart_sb.update_rbr_data(rdata);
		end

		phase.drop_objection(this);
	endtask

endclass
