interface uart_if();

  logic tx;
  logic rx;
	logic interrupt;
  
endinterface
